module fs_with_d38_tb();
reg a,b,c;
wire diff,borrow;
integer i,handle1;
fs_with_d38 dut (a,b,c,diff,borrow);
task initialize;
{a,b,c} = 3'b0;
endtask
task inputs(input[2:0]k);
begin
{a,b,c} = k;
#10;
end
endtask
initial begin
initialize;
for(i = 0; i<8; i= i+1) begin
inputs(i);
#10;
end
$fclose(handle1);
end
initial 
handle1 = $fopen("file1.txt");
initial
$fmonitor(handle1,$time, " inputs = %b %b %b ,outputs = %b %b",a,b,c,diff,borrow);
initial 
#350 $finish();
endmodule