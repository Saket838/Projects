module rst_logic(input b,c,output y);
assign y = ~(b | c);
endmodule
