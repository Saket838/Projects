module comp (a,b,greater,equal,less);
input[1:0] a,b;
output greater,equal,less;
assign greater = a[0] & ~b[1] & ~b[0] | a[1] & ~b[1] | a[1] & a[0] & ~b[0];
assign equal = ~{a[0] ^ b[0]} & ~{a[1] ^ b[1]};
assign less = ~a[1] & ~a[0] & b[0] | ~a[0] & b[1] & b[0] | ~a[1] & b[1];
endmodule
