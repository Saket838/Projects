module cla(a,b,cin,s,cout);
input[3:0] a,b;
input cin;
output [3:0] s;
output cout;
wire [3:0]c,g,p;
assign g = a & b;
assign p = a ^ b;
assign c[0] = cin;
assign c[1] = g[0] | (p[0] & c[0]);
assign c[2] = g[1] | (p[1] & g[0]) | (p[1] & p[0] & c[0]);
assign c[3] = g[2] | (p[2] & g[1]) | (p[2] & p[1] & g[0]) | (p[2] & p[1] & p[0] & c[0]);
assign cout = g[3] | (p[3] & g[2]) | (p[3] & p[2] & p[1] & g[0]) | (p[3] & p[2] & p[1] & p[0] & c[0]);
fa f1 (a[0],b[0],c[0],s[0],c[1]);
fa f2 (a[1],b[1],c[1],s[1],c[2]);
fa f3 (a[2],b[2],c[2],s[2],c[3]);
fa f4 (a[3],b[3],c[3],s[3],cout);
endmodule
