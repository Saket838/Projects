module d_ff_tb();
reg d,clk,rst;
wire q,qbar;
d_ff dut (d,clk,rst,q,qbar);
initial begin
clk = 1'b0;
forever 
#5 clk = ~clk;
end
task initialize;
begin
d = 1'b0;
rst = 1'b1;
end
endtask
task rst_dut;
begin
@ (negedge clk)
rst = 1'b1;
@ (negedge clk)
rst = 1'b0;
end
endtask
task inputs(input k);
begin
@ (negedge clk)
d = k;
end
endtask
initial begin
initialize;
rst_dut;
inputs(1'b1);
inputs(1'b0);
inputs(1'b1);
rst_dut;
end
initial #200 $finish();
endmodule
